module day_01_core (
	input wire clk,
	input wire rst,
	output reg [31:0] result,
	output reg done
);

`include "day_01_input.v"
	reg [6:0] current_position;
	reg [12:0] num_zeros;
	reg [12:0] index;

	wire [6:0] next_position;

	always @(posedge clk) begin
		if (rst) begin
			// reset to initial values
			current_position <= 50;
			num_zeros <= 0;
			index <= 0; 
			done <= 0;
			result <= 0;
		end else begin
			// normal operation
			if (index == NUM_ROTATIONS) begin
				// we're done
				done <= 1;
				result <= num_zeros;
			end else begin
				// process next rotation
				current_position <= next_position;
				if (next_position == 0) begin
					num_zeros <= num_zeros + 1;	
					end
					index <= index + 1;
				end
		end
	end

	wire direction = rotations[index][7];
	wire [6:0] distance = rotations[index][6:0]; 

	assign next_position = (direction == 0) ? ((distance > current_position) ? (100 + current_position - distance) : (current_position - distance))
											: (((current_position + distance) >= 100) ? (current_position + distance - 100) : (current_position + distance));
											
											
endmodule